// Automatically generated Verilog-2001
module Top_topEntity(input_0_0
                    ,input_0_1
                    ,// clock
                    system1000
                    ,// asynchronous reset: active low
                    system1000_rstn
                    ,output_0_0
                    ,output_0_1_0
                    ,output_0_1_1
                    ,output_0_1_2
                    ,output_0_1_3
                    ,output_0_1_4
                    ,output_0_1_5
                    ,output_0_1_6
                    ,output_0_1_7
                    ,output_0_1_8
                    ,output_0_1_9
                    ,output_0_1_10
                    ,output_0_1_11
                    ,output_0_1_12
                    ,output_0_1_13
                    ,output_0_1_14
                    ,output_0_1_15
                    ,output_0_1_16
                    ,output_0_1_17
                    ,output_0_1_18
                    ,output_0_1_19
                    ,output_0_1_20
                    ,output_0_1_21
                    ,output_0_1_22
                    ,output_0_1_23
                    ,output_0_1_24
                    ,output_0_1_25
                    ,output_0_1_26
                    ,output_0_1_27
                    ,output_0_1_28
                    ,output_0_1_29);
  input [0:0] input_0_0;
  input [0:0] input_0_1;
  input system1000;
  input system1000_rstn;
  output [0:0] output_0_0;
  output [3:0] output_0_1_0;
  output [3:0] output_0_1_1;
  output [3:0] output_0_1_2;
  output [3:0] output_0_1_3;
  output [3:0] output_0_1_4;
  output [3:0] output_0_1_5;
  output [3:0] output_0_1_6;
  output [3:0] output_0_1_7;
  output [3:0] output_0_1_8;
  output [3:0] output_0_1_9;
  output [3:0] output_0_1_10;
  output [3:0] output_0_1_11;
  output [3:0] output_0_1_12;
  output [3:0] output_0_1_13;
  output [3:0] output_0_1_14;
  output [3:0] output_0_1_15;
  output [3:0] output_0_1_16;
  output [3:0] output_0_1_17;
  output [3:0] output_0_1_18;
  output [3:0] output_0_1_19;
  output [3:0] output_0_1_20;
  output [3:0] output_0_1_21;
  output [3:0] output_0_1_22;
  output [3:0] output_0_1_23;
  output [3:0] output_0_1_24;
  output [3:0] output_0_1_25;
  output [3:0] output_0_1_26;
  output [3:0] output_0_1_27;
  output [3:0] output_0_1_28;
  output [3:0] output_0_1_29;
  wire [1:0] input_0;
  wire [120:0] output_0;
  wire [119:0] output_0_1;
  assign input_0 = {input_0_0
                   ,input_0_1};
  
  Top_topEntity_0 Top_topEntity_0_inst
  (.arg (input_0)
  ,.system1000 (system1000)
  ,.system1000_rstn (system1000_rstn)
  ,.result (output_0));
  
  assign output_0_0 = output_0[120:120];
  
  assign output_0_1 = output_0[119:0];
  
  assign output_0_1_0 = output_0_1[119:116];
  
  assign output_0_1_1 = output_0_1[115:112];
  
  assign output_0_1_2 = output_0_1[111:108];
  
  assign output_0_1_3 = output_0_1[107:104];
  
  assign output_0_1_4 = output_0_1[103:100];
  
  assign output_0_1_5 = output_0_1[99:96];
  
  assign output_0_1_6 = output_0_1[95:92];
  
  assign output_0_1_7 = output_0_1[91:88];
  
  assign output_0_1_8 = output_0_1[87:84];
  
  assign output_0_1_9 = output_0_1[83:80];
  
  assign output_0_1_10 = output_0_1[79:76];
  
  assign output_0_1_11 = output_0_1[75:72];
  
  assign output_0_1_12 = output_0_1[71:68];
  
  assign output_0_1_13 = output_0_1[67:64];
  
  assign output_0_1_14 = output_0_1[63:60];
  
  assign output_0_1_15 = output_0_1[59:56];
  
  assign output_0_1_16 = output_0_1[55:52];
  
  assign output_0_1_17 = output_0_1[51:48];
  
  assign output_0_1_18 = output_0_1[47:44];
  
  assign output_0_1_19 = output_0_1[43:40];
  
  assign output_0_1_20 = output_0_1[39:36];
  
  assign output_0_1_21 = output_0_1[35:32];
  
  assign output_0_1_22 = output_0_1[31:28];
  
  assign output_0_1_23 = output_0_1[27:24];
  
  assign output_0_1_24 = output_0_1[23:20];
  
  assign output_0_1_25 = output_0_1[19:16];
  
  assign output_0_1_26 = output_0_1[15:12];
  
  assign output_0_1_27 = output_0_1[11:8];
  
  assign output_0_1_28 = output_0_1[7:4];
  
  assign output_0_1_29 = output_0_1[3:0];
endmodule
